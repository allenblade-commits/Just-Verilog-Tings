// This module outputs a constant logic LOW (0).
module top_module(output zero);
    
    // Assigning the output 'zero' a constant value of 1'b0 (binary 0).
    assign zero = 1'b0;
    
endmodule
